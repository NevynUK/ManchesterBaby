/************************************************
*  Manchester Baby in System Verilog            *
*  Richard Leivers - July 2009                  *
*                                               *
*  NIGHT PROGRAM MEMORY FILE                    *
*  Automatically generated from NIGHT.SNP       *
*                                               *
************************************************/

module progNIGHT (
    output reg signed [31:0] prog [0:31]
    );

    reverser r0 (.in(32'b00000110101001000100000100000100),.out(prog[0][31:0]));
    reverser r1 (.in(32'b10011011111100100010000010001000),.out(prog[1][31:0]));
    reverser r2 (.in(32'b10000010000101101000100001010000),.out(prog[2][31:0]));
    reverser r3 (.in(32'b00000010000100110100001001100000),.out(prog[3][31:0]));
    reverser r4 (.in(32'b11101011111100011010101010010100),.out(prog[4][31:0]));
    reverser r5 (.in(32'b10000000110000010001000010101001),.out(prog[5][31:0]));
    reverser r6 (.in(32'b10000001111000010000100100001100),.out(prog[6][31:0]));
    reverser r7 (.in(32'b10000001111000010000011000000010),.out(prog[7][31:0]));
    reverser r8 (.in(32'b10011000000001101000011001000001),.out(prog[8][31:0]));
    reverser r9 (.in(32'b10101001111000100100100100000010),.out(prog[9][31:0]));
    reverser r10 (.in(32'b00000001111000110011010010000100),.out(prog[10][31:0]));
    reverser r11 (.in(32'b01101001111000010011000001001000),.out(prog[11][31:0]));
    reverser r12 (.in(32'b11101001111000010100100000110000),.out(prog[12][31:0]));
    reverser r13 (.in(32'b10101000110001101000010000110000),.out(prog[13][31:0]));
    reverser r14 (.in(32'b10100001111000010000001001001000),.out(prog[14][31:0]));
    reverser r15 (.in(32'b00010011111101100000000110000100),.out(prog[15][31:0]));
    reverser r16 (.in(32'b00000111111110010000000010000010),.out(prog[16][31:0]));
    reverser r17 (.in(32'b10000011111101101111111111111111),.out(prog[17][31:0]));
    reverser r18 (.in(32'b10101001111000100110011001100110),.out(prog[18][31:0]));
    reverser r19 (.in(32'b10101000110001101111111111111111),.out(prog[19][31:0]));
    reverser r20 (.in(32'b00011000110000001111111111111111),.out(prog[20][31:0]));
    reverser r21 (.in(32'b01100000000000000000000000000000),.out(prog[21][31:0]));
    reverser r22 (.in(32'b11100000000000000000000000000000),.out(prog[22][31:0]));
    reverser r23 (.in(32'b11111111111111111111111111111111),.out(prog[23][31:0]));
    reverser r24 (.in(32'b00000000000000000000000000000000),.out(prog[24][31:0]));
    reverser r25 (.in(32'b00000000000000011111000000100000),.out(prog[25][31:0]));
    reverser r26 (.in(32'b00000000000000100000100001010000),.out(prog[26][31:0]));
    reverser r27 (.in(32'b00000000000000100010100000100000),.out(prog[27][31:0]));
    reverser r28 (.in(32'b00000001111110100000100000111000),.out(prog[28][31:0]));
    reverser r29 (.in(32'b00000010000000011111000000100000),.out(prog[29][31:0]));
    reverser r30 (.in(32'b00011110011110001000000000100000),.out(prog[30][31:0]));
    reverser r31 (.in(32'b00111111111111111110000001010000),.out(prog[31][31:0]));

endmodule
