/************************************************ 	
 *	Manchester Baby in System Verilog  			*
 * 	Richard Leivers - July 2009        			*
 * 												*
 *	PARABOLA PROGRAM MEMORY FILE				*
 *  Automatically generated from PARABOLA.SNP	*
 *												*
 ************************************************/
 
 module progPARABOLA (
	output reg signed [31:0] prog [0:31]
	);
	
	reverser r0 (.in(32'b00000000000000000000000000000000),.out(prog[0][31:0]));
	reverser r1 (.in(32'b10111000000000100000000000000000),.out(prog[1][31:0]));	
	reverser r2 (.in(32'b10111000000000010000000000000000),.out(prog[2][31:0]));	
	reverser r3 (.in(32'b10111000000001100000000000000000),.out(prog[3][31:0]));	
	reverser r4 (.in(32'b00000000000000110000000000000000),.out(prog[4][31:0]));	
	reverser r5 (.in(32'b00000000000001110000000000000000),.out(prog[5][31:0]));
	reverser r6 (.in(32'b10111000000000100000000000000000),.out(prog[6][31:0]));
	reverser r7 (.in(32'b10111000000001100000000000000000),.out(prog[7][31:0]));
	reverser r8 (.in(32'b01101000000000100000000000000000),.out(prog[8][31:0]));
	reverser r9 (.in(32'b10111000000000010000000000000000),.out(prog[9][31:0]));
	reverser r10 (.in(32'b01111000000001100000000000000000),.out(prog[10][31:0]));
	reverser r11 (.in(32'b01111000000000100000000000000000),.out(prog[11][31:0]));
	reverser r12 (.in(32'b01101000000001100000000000000000),.out(prog[12][31:0]));
	reverser r13 (.in(32'b00010000000000100000000000000000),.out(prog[13][31:0]));
	reverser r14 (.in(32'b00111000000000010000000000000000),.out(prog[14][31:0]));	
	reverser r15 (.in(32'b01111000000001100000000000000000),.out(prog[15][31:0]));	
	reverser r16 (.in(32'b01111000000000100000000000000000),.out(prog[16][31:0]));
	reverser r17 (.in(32'b00010000000001100000000000000000),.out(prog[17][31:0]));
	reverser r18 (.in(32'b11011000000000010000000000000000),.out(prog[18][31:0]));
	reverser r19 (.in(32'b00110000000001100000000000000000),.out(prog[19][31:0]));
	reverser r20 (.in(32'b00111000000000100000000000000000),.out(prog[20][31:0]));
	reverser r21 (.in(32'b01011000000000010000000000000000),.out(prog[21][31:0]));
	reverser r22 (.in(32'b00111000000001100000000000000000),.out(prog[22][31:0]));
	reverser r23 (.in(32'b00111000000000100000000000000000),.out(prog[23][31:0]));
	reverser r24 (.in(32'b00111000000001100000000000000000),.out(prog[24][31:0]));
	reverser r25 (.in(32'b11111000000000000000000000000000),.out(prog[25][31:0]));	
	reverser r26 (.in(32'b10000000000000000000000000000000),.out(prog[26][31:0]));
	reverser r27 (.in(32'b00000000000001111111111111111111),.out(prog[27][31:0]));
	reverser r28 (.in(32'b01011111111111111111111111111111),.out(prog[28][31:0]));	
	reverser r29 (.in(32'b00000000000000000100000000000000),.out(prog[29][31:0]));	
	reverser r30 (.in(32'b00000000000000000000000000000000),.out(prog[30][31:0]));	
	reverser r31 (.in(32'b00000000000000000000000000000000),.out(prog[31][31:0]));

endmodule
